module PPGenerator( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input         io_in_input_sign, // @[:@6.4]
  input  [7:0]  io_in_input_exponent, // @[:@6.4]
  input  [22:0] io_in_input_mantissa, // @[:@6.4]
  input  [2:0]  io_in_weight_grps_0, // @[:@6.4]
  input  [2:0]  io_in_weight_grps_1, // @[:@6.4]
  input  [7:0]  io_in_weight_exponent, // @[:@6.4]
  output [12:0] io_out_pp_1, // @[:@6.4]
  output [12:0] io_out_pp_2, // @[:@6.4]
  output [8:0]  io_out_exponent // @[:@6.4]
);
  wire [1:0] _T_47; // @[PPGenerator.scala 24:38:@10.4]
  wire  _T_49; // @[PPGenerator.scala 24:44:@11.4]
  wire [2:0] _T_52; // @[PPGenerator.scala 24:97:@12.4]
  wire [3:0] _T_53; // @[Cat.scala 30:58:@13.4]
  wire [6:0] _GEN_0; // @[PPGenerator.scala 24:106:@15.4]
  wire [6:0] _T_55; // @[PPGenerator.scala 24:106:@15.4]
  wire [9:0] _GEN_1; // @[PPGenerator.scala 24:135:@16.4]
  wire [9:0] _T_56; // @[PPGenerator.scala 24:135:@16.4]
  wire [9:0] _T_57; // @[PPGenerator.scala 24:17:@17.4]
  wire [1:0] _T_58; // @[PPGenerator.scala 25:38:@19.4]
  wire  _T_60; // @[PPGenerator.scala 25:44:@20.4]
  wire [6:0] _T_66; // @[PPGenerator.scala 25:106:@24.4]
  wire [6:0] _T_67; // @[PPGenerator.scala 25:17:@25.4]
  wire  _T_68; // @[PPGenerator.scala 27:61:@27.4]
  wire  _T_69; // @[PPGenerator.scala 27:39:@28.4]
  wire [8:0] pp1_tmp; // @[PPGenerator.scala 21:21:@8.4 PPGenerator.scala 24:11:@18.4]
  wire [9:0] _T_70; // @[Cat.scala 30:58:@29.4]
  wire [8:0] pp2_tmp; // @[PPGenerator.scala 22:21:@9.4 PPGenerator.scala 25:11:@26.4]
  wire [9:0] _T_73; // @[Cat.scala 30:58:@33.4]
  wire [8:0] _T_74; // @[PPGenerator.scala 29:43:@35.4]
  wire [7:0] _T_75; // @[PPGenerator.scala 29:43:@36.4]
  assign _T_47 = io_in_weight_grps_1[1:0]; // @[PPGenerator.scala 24:38:@10.4]
  assign _T_49 = _T_47 == 2'h3; // @[PPGenerator.scala 24:44:@11.4]
  assign _T_52 = io_in_input_mantissa[22:20]; // @[PPGenerator.scala 24:97:@12.4]
  assign _T_53 = {1'h1,_T_52}; // @[Cat.scala 30:58:@13.4]
  assign _GEN_0 = {{3'd0}, _T_53}; // @[PPGenerator.scala 24:106:@15.4]
  assign _T_55 = _GEN_0 << _T_47; // @[PPGenerator.scala 24:106:@15.4]
  assign _GEN_1 = {{3'd0}, _T_55}; // @[PPGenerator.scala 24:135:@16.4]
  assign _T_56 = _GEN_1 << 3; // @[PPGenerator.scala 24:135:@16.4]
  assign _T_57 = _T_49 ? 10'h0 : _T_56; // @[PPGenerator.scala 24:17:@17.4]
  assign _T_58 = io_in_weight_grps_0[1:0]; // @[PPGenerator.scala 25:38:@19.4]
  assign _T_60 = _T_58 == 2'h3; // @[PPGenerator.scala 25:44:@20.4]
  assign _T_66 = _GEN_0 << _T_58; // @[PPGenerator.scala 25:106:@24.4]
  assign _T_67 = _T_60 ? 7'h0 : _T_66; // @[PPGenerator.scala 25:17:@25.4]
  assign _T_68 = io_in_weight_grps_1[2]; // @[PPGenerator.scala 27:61:@27.4]
  assign _T_69 = io_in_input_sign ^ _T_68; // @[PPGenerator.scala 27:39:@28.4]
  assign pp1_tmp = _T_57[8:0]; // @[PPGenerator.scala 21:21:@8.4 PPGenerator.scala 24:11:@18.4]
  assign _T_70 = {_T_69,pp1_tmp}; // @[Cat.scala 30:58:@29.4]
  assign pp2_tmp = {{2'd0}, _T_67}; // @[PPGenerator.scala 22:21:@9.4 PPGenerator.scala 25:11:@26.4]
  assign _T_73 = {_T_69,pp2_tmp}; // @[Cat.scala 30:58:@33.4]
  assign _T_74 = io_in_input_exponent + io_in_weight_exponent; // @[PPGenerator.scala 29:43:@35.4]
  assign _T_75 = _T_74[7:0]; // @[PPGenerator.scala 29:43:@36.4]
  assign io_out_pp_1 = {{3'd0}, _T_70}; // @[PPGenerator.scala 27:15:@30.4]
  assign io_out_pp_2 = {{3'd0}, _T_73}; // @[PPGenerator.scala 28:15:@34.4]
  assign io_out_exponent = {{1'd0}, _T_75}; // @[PPGenerator.scala 29:19:@37.4]
endmodule
