module SignAdder( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [17:0] io_in, // @[:@6.4]
  output [5:0]  io_out // @[:@6.4]
);
  wire  _T_40; // @[Signadder.scala 15:22:@12.4]
  wire  _T_41; // @[Signadder.scala 15:35:@13.4]
  wire [1:0] _T_42; // @[Signadder.scala 15:28:@14.4]
  wire  _T_43; // @[Signadder.scala 15:28:@15.4]
  wire  _T_44; // @[Signadder.scala 15:22:@17.4]
  wire  _T_45; // @[Signadder.scala 15:35:@18.4]
  wire [1:0] _T_46; // @[Signadder.scala 15:28:@19.4]
  wire  _T_47; // @[Signadder.scala 15:28:@20.4]
  wire  _T_48; // @[Signadder.scala 15:22:@22.4]
  wire  _T_49; // @[Signadder.scala 15:35:@23.4]
  wire [1:0] _T_50; // @[Signadder.scala 15:28:@24.4]
  wire  _T_51; // @[Signadder.scala 15:28:@25.4]
  wire  _T_52; // @[Signadder.scala 15:22:@27.4]
  wire  _T_53; // @[Signadder.scala 15:35:@28.4]
  wire [1:0] _T_54; // @[Signadder.scala 15:28:@29.4]
  wire  _T_55; // @[Signadder.scala 15:28:@30.4]
  wire  _T_56; // @[Signadder.scala 15:22:@32.4]
  wire  _T_57; // @[Signadder.scala 15:35:@33.4]
  wire [1:0] _T_58; // @[Signadder.scala 15:28:@34.4]
  wire  _T_59; // @[Signadder.scala 15:28:@35.4]
  wire  _T_60; // @[Signadder.scala 15:22:@37.4]
  wire  _T_61; // @[Signadder.scala 15:35:@38.4]
  wire [1:0] _T_62; // @[Signadder.scala 15:28:@39.4]
  wire  _T_63; // @[Signadder.scala 15:28:@40.4]
  wire  _T_64; // @[Signadder.scala 15:22:@42.4]
  wire  _T_65; // @[Signadder.scala 15:35:@43.4]
  wire [1:0] _T_66; // @[Signadder.scala 15:28:@44.4]
  wire  _T_67; // @[Signadder.scala 15:28:@45.4]
  wire  _T_68; // @[Signadder.scala 15:22:@47.4]
  wire  _T_69; // @[Signadder.scala 15:35:@48.4]
  wire [1:0] _T_70; // @[Signadder.scala 15:28:@49.4]
  wire  _T_71; // @[Signadder.scala 15:28:@50.4]
  wire  _T_72; // @[Signadder.scala 15:22:@52.4]
  wire  _T_73; // @[Signadder.scala 15:35:@53.4]
  wire [1:0] _T_74; // @[Signadder.scala 15:28:@54.4]
  wire  _T_75; // @[Signadder.scala 15:28:@55.4]
  wire [1:0] tmp_1_0; // @[Signadder.scala 10:19:@8.4 Signadder.scala 15:14:@16.4]
  wire [1:0] tmp_1_1; // @[Signadder.scala 10:19:@8.4 Signadder.scala 15:14:@21.4]
  wire [2:0] _T_76; // @[Signadder.scala 18:28:@57.4]
  wire [1:0] _T_77; // @[Signadder.scala 18:28:@58.4]
  wire [1:0] tmp_1_2; // @[Signadder.scala 10:19:@8.4 Signadder.scala 15:14:@26.4]
  wire [1:0] tmp_1_3; // @[Signadder.scala 10:19:@8.4 Signadder.scala 15:14:@31.4]
  wire [2:0] _T_78; // @[Signadder.scala 18:28:@60.4]
  wire [1:0] _T_79; // @[Signadder.scala 18:28:@61.4]
  wire [1:0] tmp_1_4; // @[Signadder.scala 10:19:@8.4 Signadder.scala 15:14:@36.4]
  wire [1:0] tmp_1_5; // @[Signadder.scala 10:19:@8.4 Signadder.scala 15:14:@41.4]
  wire [2:0] _T_80; // @[Signadder.scala 18:28:@63.4]
  wire [1:0] _T_81; // @[Signadder.scala 18:28:@64.4]
  wire [1:0] tmp_1_6; // @[Signadder.scala 10:19:@8.4 Signadder.scala 15:14:@46.4]
  wire [1:0] tmp_1_7; // @[Signadder.scala 10:19:@8.4 Signadder.scala 15:14:@51.4]
  wire [2:0] _T_82; // @[Signadder.scala 18:28:@66.4]
  wire [1:0] _T_83; // @[Signadder.scala 18:28:@67.4]
  wire [2:0] tmp_2_0; // @[Signadder.scala 11:19:@9.4 Signadder.scala 18:14:@59.4]
  wire [2:0] tmp_2_1; // @[Signadder.scala 11:19:@9.4 Signadder.scala 18:14:@62.4]
  wire [3:0] _T_84; // @[Signadder.scala 21:28:@69.4]
  wire [2:0] _T_85; // @[Signadder.scala 21:28:@70.4]
  wire [2:0] tmp_2_2; // @[Signadder.scala 11:19:@9.4 Signadder.scala 18:14:@65.4]
  wire [2:0] tmp_2_3; // @[Signadder.scala 11:19:@9.4 Signadder.scala 18:14:@68.4]
  wire [3:0] _T_86; // @[Signadder.scala 21:28:@72.4]
  wire [2:0] _T_87; // @[Signadder.scala 21:28:@73.4]
  wire [3:0] tmp_3_0; // @[Signadder.scala 12:19:@10.4 Signadder.scala 21:14:@71.4]
  wire [3:0] tmp_3_1; // @[Signadder.scala 12:19:@10.4 Signadder.scala 21:14:@74.4]
  wire [4:0] _T_88; // @[Signadder.scala 23:21:@75.4]
  wire [3:0] _T_89; // @[Signadder.scala 23:21:@76.4]
  wire [4:0] tmp_4; // @[Signadder.scala 13:19:@11.4 Signadder.scala 23:9:@77.4]
  wire [1:0] tmp_1_8; // @[Signadder.scala 10:19:@8.4 Signadder.scala 15:14:@56.4]
  wire [4:0] _GEN_0; // @[Signadder.scala 24:20:@78.4]
  wire [5:0] _T_90; // @[Signadder.scala 24:20:@78.4]
  wire [5:0] _T_91; // @[Signadder.scala 24:13:@79.4]
  wire [6:0] _T_93; // @[Signadder.scala 24:32:@80.4]
  assign _T_40 = io_in[0]; // @[Signadder.scala 15:22:@12.4]
  assign _T_41 = io_in[1]; // @[Signadder.scala 15:35:@13.4]
  assign _T_42 = _T_40 + _T_41; // @[Signadder.scala 15:28:@14.4]
  assign _T_43 = _T_42[0:0]; // @[Signadder.scala 15:28:@15.4]
  assign _T_44 = io_in[2]; // @[Signadder.scala 15:22:@17.4]
  assign _T_45 = io_in[3]; // @[Signadder.scala 15:35:@18.4]
  assign _T_46 = _T_44 + _T_45; // @[Signadder.scala 15:28:@19.4]
  assign _T_47 = _T_46[0:0]; // @[Signadder.scala 15:28:@20.4]
  assign _T_48 = io_in[4]; // @[Signadder.scala 15:22:@22.4]
  assign _T_49 = io_in[5]; // @[Signadder.scala 15:35:@23.4]
  assign _T_50 = _T_48 + _T_49; // @[Signadder.scala 15:28:@24.4]
  assign _T_51 = _T_50[0:0]; // @[Signadder.scala 15:28:@25.4]
  assign _T_52 = io_in[6]; // @[Signadder.scala 15:22:@27.4]
  assign _T_53 = io_in[7]; // @[Signadder.scala 15:35:@28.4]
  assign _T_54 = _T_52 + _T_53; // @[Signadder.scala 15:28:@29.4]
  assign _T_55 = _T_54[0:0]; // @[Signadder.scala 15:28:@30.4]
  assign _T_56 = io_in[8]; // @[Signadder.scala 15:22:@32.4]
  assign _T_57 = io_in[9]; // @[Signadder.scala 15:35:@33.4]
  assign _T_58 = _T_56 + _T_57; // @[Signadder.scala 15:28:@34.4]
  assign _T_59 = _T_58[0:0]; // @[Signadder.scala 15:28:@35.4]
  assign _T_60 = io_in[10]; // @[Signadder.scala 15:22:@37.4]
  assign _T_61 = io_in[11]; // @[Signadder.scala 15:35:@38.4]
  assign _T_62 = _T_60 + _T_61; // @[Signadder.scala 15:28:@39.4]
  assign _T_63 = _T_62[0:0]; // @[Signadder.scala 15:28:@40.4]
  assign _T_64 = io_in[12]; // @[Signadder.scala 15:22:@42.4]
  assign _T_65 = io_in[13]; // @[Signadder.scala 15:35:@43.4]
  assign _T_66 = _T_64 + _T_65; // @[Signadder.scala 15:28:@44.4]
  assign _T_67 = _T_66[0:0]; // @[Signadder.scala 15:28:@45.4]
  assign _T_68 = io_in[14]; // @[Signadder.scala 15:22:@47.4]
  assign _T_69 = io_in[15]; // @[Signadder.scala 15:35:@48.4]
  assign _T_70 = _T_68 + _T_69; // @[Signadder.scala 15:28:@49.4]
  assign _T_71 = _T_70[0:0]; // @[Signadder.scala 15:28:@50.4]
  assign _T_72 = io_in[16]; // @[Signadder.scala 15:22:@52.4]
  assign _T_73 = io_in[17]; // @[Signadder.scala 15:35:@53.4]
  assign _T_74 = _T_72 + _T_73; // @[Signadder.scala 15:28:@54.4]
  assign _T_75 = _T_74[0:0]; // @[Signadder.scala 15:28:@55.4]
  assign tmp_1_0 = {{1'd0}, _T_43}; // @[Signadder.scala 10:19:@8.4 Signadder.scala 15:14:@16.4]
  assign tmp_1_1 = {{1'd0}, _T_47}; // @[Signadder.scala 10:19:@8.4 Signadder.scala 15:14:@21.4]
  assign _T_76 = tmp_1_0 + tmp_1_1; // @[Signadder.scala 18:28:@57.4]
  assign _T_77 = _T_76[1:0]; // @[Signadder.scala 18:28:@58.4]
  assign tmp_1_2 = {{1'd0}, _T_51}; // @[Signadder.scala 10:19:@8.4 Signadder.scala 15:14:@26.4]
  assign tmp_1_3 = {{1'd0}, _T_55}; // @[Signadder.scala 10:19:@8.4 Signadder.scala 15:14:@31.4]
  assign _T_78 = tmp_1_2 + tmp_1_3; // @[Signadder.scala 18:28:@60.4]
  assign _T_79 = _T_78[1:0]; // @[Signadder.scala 18:28:@61.4]
  assign tmp_1_4 = {{1'd0}, _T_59}; // @[Signadder.scala 10:19:@8.4 Signadder.scala 15:14:@36.4]
  assign tmp_1_5 = {{1'd0}, _T_63}; // @[Signadder.scala 10:19:@8.4 Signadder.scala 15:14:@41.4]
  assign _T_80 = tmp_1_4 + tmp_1_5; // @[Signadder.scala 18:28:@63.4]
  assign _T_81 = _T_80[1:0]; // @[Signadder.scala 18:28:@64.4]
  assign tmp_1_6 = {{1'd0}, _T_67}; // @[Signadder.scala 10:19:@8.4 Signadder.scala 15:14:@46.4]
  assign tmp_1_7 = {{1'd0}, _T_71}; // @[Signadder.scala 10:19:@8.4 Signadder.scala 15:14:@51.4]
  assign _T_82 = tmp_1_6 + tmp_1_7; // @[Signadder.scala 18:28:@66.4]
  assign _T_83 = _T_82[1:0]; // @[Signadder.scala 18:28:@67.4]
  assign tmp_2_0 = {{1'd0}, _T_77}; // @[Signadder.scala 11:19:@9.4 Signadder.scala 18:14:@59.4]
  assign tmp_2_1 = {{1'd0}, _T_79}; // @[Signadder.scala 11:19:@9.4 Signadder.scala 18:14:@62.4]
  assign _T_84 = tmp_2_0 + tmp_2_1; // @[Signadder.scala 21:28:@69.4]
  assign _T_85 = _T_84[2:0]; // @[Signadder.scala 21:28:@70.4]
  assign tmp_2_2 = {{1'd0}, _T_81}; // @[Signadder.scala 11:19:@9.4 Signadder.scala 18:14:@65.4]
  assign tmp_2_3 = {{1'd0}, _T_83}; // @[Signadder.scala 11:19:@9.4 Signadder.scala 18:14:@68.4]
  assign _T_86 = tmp_2_2 + tmp_2_3; // @[Signadder.scala 21:28:@72.4]
  assign _T_87 = _T_86[2:0]; // @[Signadder.scala 21:28:@73.4]
  assign tmp_3_0 = {{1'd0}, _T_85}; // @[Signadder.scala 12:19:@10.4 Signadder.scala 21:14:@71.4]
  assign tmp_3_1 = {{1'd0}, _T_87}; // @[Signadder.scala 12:19:@10.4 Signadder.scala 21:14:@74.4]
  assign _T_88 = tmp_3_0 + tmp_3_1; // @[Signadder.scala 23:21:@75.4]
  assign _T_89 = _T_88[3:0]; // @[Signadder.scala 23:21:@76.4]
  assign tmp_4 = {{1'd0}, _T_89}; // @[Signadder.scala 13:19:@11.4 Signadder.scala 23:9:@77.4]
  assign tmp_1_8 = {{1'd0}, _T_75}; // @[Signadder.scala 10:19:@8.4 Signadder.scala 15:14:@56.4]
  assign _GEN_0 = {{3'd0}, tmp_1_8}; // @[Signadder.scala 24:20:@78.4]
  assign _T_90 = tmp_4 + _GEN_0; // @[Signadder.scala 24:20:@78.4]
  assign _T_91 = ~ _T_90; // @[Signadder.scala 24:13:@79.4]
  assign _T_93 = _T_91 + 6'h1; // @[Signadder.scala 24:32:@80.4]
  assign io_out = _T_93[5:0]; // @[Signadder.scala 24:10:@82.4]
endmodule
